interface pds_if(input clk);
	logic req;
	logic fault;
	logic gnt;
endinterface