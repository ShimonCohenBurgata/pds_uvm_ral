

package pds_env_pkg;
	import uvm_pkg::*;
	`include "uvm_macros.svh"

	import apb_agent_pkg::*;
	import pds_agent_pkg::*;
	import pds_reg_pkg::*;

	`include "pds_env_config.svh"
	`include "reg_env.svh"
	`include "pds_scoreboard.svh"
	`include "pds_env.svh"

endpackage:pds_env_pkg