

package pds_test_lib_pkg;
	
	import uvm_pkg::*;
	`include "uvm_macros.svh"
	
	import pds_env_pkg::*;
	import apb_agent_pkg::*;
	import pds_agent_pkg::*;
	import apb_bus_sequence_lib_pkg::*;
	import pds_reg_pkg::*;
	
		
	`include "pds_test_base.svh"
	`include "pds_simple_test.svh"
endpackage:pds_test_lib_pkg