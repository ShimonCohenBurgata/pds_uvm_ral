

module hvl_top;
	import uvm_pkg::*;
	import pds_test_lib_pkg::*;
	
	initial begin
		run_test("pds_simple_test");
	end
endmodule:hvl_top